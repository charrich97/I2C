package wb_pkg;
	import utility_pkg::*;
	import ncsu_pkg::*;
	`include "../../../ncsu_pkg/ncsu_macros.svh"
  `include "UVM/wb_configuration.svh"
  `include "UVM/wb_transaction.svh"
  `include "UVM/wb_driver.svh"
  `include "UVM/wb_monitor.svh"
	`include "UVM/wb_sequence.svh"
	`include "UVM/wb_coverage_sequence.svh"
  `include "UVM/wb_random_sequence.svh"
  `include "UVM/wb_agent.svh"
endpackage
