package i2c_pkg;
  import utility_pkg::*;
  import ncsu_pkg::*;
  `include "../../../ncsu_pkg/ncsu_macros.svh"
  `include "UVM/i2c_configuration.svh"
  `include "UVM/i2c_transaction.svh"
  `include "UVM/i2c_driver.svh"
  `include "UVM/i2c_monitor.svh"
  `include "UVM/i2c_sequence.svh"
  `include "UVM/i2c_coverage_sequence.svh"
  `include "UVM/i2c_random_sequence.svh"
  `include "UVM/i2c_agent.svh"
endpackage
