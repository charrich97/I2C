package i2cmb_env_pkg;
	import ncsu_pkg::*;
	import utility_pkg::*;
	import wb_pkg::*;
	import i2c_pkg::*;
	`include "../../../ncsu_pkg/ncsu_macros.svh"
  `include "UVM/i2cmb_env_configuration.svh"
  `include "UVM/i2cmb_generator.svh"
  `include "UVM/i2cmb_predictor.svh"
  `include "UVM/i2cmb_scoreboard.svh"
  `include "UVM/i2cmb_coverage.svh"
  `include "UVM/i2cmb_environment.svh"
  `include "UVM/i2cmb_test.svh"
endpackage //i2cmb_env_pkg
